`timescale 1ns/100ps
// ============================================================
// Toy Saturnin Round - Fully Flattened (No Submodules)
// ============================================================
module APN_ANF (
    input  [31:0] state_in,
    output [31:0] state_out
);
    // ---------------------------------------------------------
    // Unpack 8 nibbles
    // ---------------------------------------------------------
    wire [3:0] x0 = state_in[31:28];
    wire [3:0] x1 = state_in[27:24];
    wire [3:0] x2 = state_in[23:20];
    wire [3:0] x3 = state_in[19:16];
    wire [3:0] x4 = state_in[15:12];
    wire [3:0] x5 = state_in[11:8];
    wire [3:0] x6 = state_in[7:4];
    wire [3:0] x7 = state_in[3:0];

    // =========================================================
    // Helper: inline APN_ANF function as a macro
    // =========================================================
    `define APN_ANF(a) { \
        ((a[0]&a[1]&a[2])^(a[0]&a[1])^(a[0]&a[2])^(a[1]&a[3])^(a[1])^(a[2])^(a[3])), \
        ((a[0]&a[2]&a[3])^(a[0]&a[2])^(a[0]&a[3])^(a[0])^(a[1]&a[2])^(a[1])^(a[2]&a[3])^(a[2])), \
        ((a[0]&a[3])^(a[0])^(a[1]&a[2]&a[3])^(a[1]&a[2])^(a[1]&a[3])^(a[1])^(a[2])), \
        ((a[0]&a[1]&a[3])^(a[0]&a[1])^(a[0]&a[2])^(a[0]&a[3])^(a[1]&a[3])^(a[2])^(a[3])) }

    // =========================================================
    // First S-box layer (8 parallel)
    // =========================================================
    wire [3:0] s1_0 = `APN_ANF(x0);
    wire [3:0] s1_1 = `APN_ANF(x1);
    wire [3:0] s1_2 = `APN_ANF(x2);
    wire [3:0] s1_3 = `APN_ANF(x3);
    wire [3:0] s1_4 = `APN_ANF(x4);
    wire [3:0] s1_5 = `APN_ANF(x5);
    wire [3:0] s1_6 = `APN_ANF(x6);
    wire [3:0] s1_7 = `APN_ANF(x7);

    // =========================================================
    // MDS Layer 1
    // =========================================================
    wire [3:0] m1_0 = s1_0 ^ s1_1 ^ s1_2 ^ s1_4 ^ s1_6;
    wire [3:0] m1_1 = s1_0 ^ s1_3 ^ s1_5 ^ s1_7;
    wire [3:0] m1_2 = s1_0 ^ s1_2 ^ s1_3 ^ s1_5;
    wire [3:0] m1_3 = s1_1 ^ s1_2 ^ s1_4 ^ s1_5;
    wire [3:0] m1_4 = s1_0 ^ s1_2 ^ s1_4 ^ s1_5 ^ s1_6;
    wire [3:0] m1_5 = s1_1 ^ s1_3 ^ s1_4 ^ s1_7;
    wire [3:0] m1_6 = s1_1 ^ s1_4 ^ s1_6 ^ s1_7;
    wire [3:0] m1_7 = s1_0 ^ s1_1 ^ s1_5 ^ s1_6;

    // =========================================================
    // Second S-box layer
    // =========================================================
    wire [3:0] s2_0 = `APN_ANF(m1_0);
    wire [3:0] s2_1 = `APN_ANF(m1_1);
    wire [3:0] s2_2 = `APN_ANF(m1_2);
    wire [3:0] s2_3 = `APN_ANF(m1_3);
    wire [3:0] s2_4 = `APN_ANF(m1_4);
    wire [3:0] s2_5 = `APN_ANF(m1_5);
    wire [3:0] s2_6 = `APN_ANF(m1_6);
    wire [3:0] s2_7 = `APN_ANF(m1_7);

    // =========================================================
    // SR_sheet (permute 4..7)
    // =========================================================
    wire [3:0] sr_0 = s2_0;
    wire [3:0] sr_1 = s2_1;
    wire [3:0] sr_2 = s2_2;
    wire [3:0] sr_3 = s2_3;
    wire [3:0] sr_4 = {s2_4[2], s2_4[3], s2_4[0], s2_4[1]};
    wire [3:0] sr_5 = {s2_5[2], s2_5[3], s2_5[0], s2_5[1]};
    wire [3:0] sr_6 = {s2_6[2], s2_6[3], s2_6[0], s2_6[1]};
    wire [3:0] sr_7 = {s2_7[2], s2_7[3], s2_7[0], s2_7[1]};

    // =========================================================
    // MDS Layer 2
    // =========================================================
    wire [3:0] m2_0 = sr_0 ^ sr_1 ^ sr_2 ^ sr_4 ^ sr_6;
    wire [3:0] m2_1 = sr_0 ^ sr_3 ^ sr_5 ^ sr_7;
    wire [3:0] m2_2 = sr_0 ^ sr_2 ^ sr_3 ^ sr_5;
    wire [3:0] m2_3 = sr_1 ^ sr_2 ^ sr_4 ^ sr_5;
    wire [3:0] m2_4 = sr_0 ^ sr_2 ^ sr_4 ^ sr_5 ^ sr_6;
    wire [3:0] m2_5 = sr_1 ^ sr_3 ^ sr_4 ^ sr_7;
    wire [3:0] m2_6 = sr_1 ^ sr_4 ^ sr_6 ^ sr_7;
    wire [3:0] m2_7 = sr_0 ^ sr_1 ^ sr_5 ^ sr_6;

    // =========================================================
    // INV_SR_sheet (same as SR_sheet)
    // =========================================================
    wire [3:0] z0 = m2_0;
    wire [3:0] z1 = m2_1;
    wire [3:0] z2 = m2_2;
    wire [3:0] z3 = m2_3;
    wire [3:0] z4 = {m2_4[2], m2_4[3], m2_4[0], m2_4[1]};
    wire [3:0] z5 = {m2_5[2], m2_5[3], m2_5[0], m2_5[1]};
    wire [3:0] z6 = {m2_6[2], m2_6[3], m2_6[0], m2_6[1]};
    wire [3:0] z7 = {m2_7[2], m2_7[3], m2_7[0], m2_7[1]};

    // =========================================================
    // Pack 8 nibbles back into 32-bit output
    // =========================================================
    assign state_out = {z0, z1, z2, z3, z4, z5, z6, z7};

endmodule
